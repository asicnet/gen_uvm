

  string seq_name = "master_init_seq";
  int    seq_var  = 0;
  string seq_mode = "nop";

  function void init_item();

  endfunction
