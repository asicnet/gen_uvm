
library IEEE;
use IEEE.std_Logic_1164.all;
use IEEE.numeric_std.all;

entity dut_top_entity is

end;

architecture rtl of dut_top_entity  is

begin

end;  
